module game(
    input system_clk, start, 
    input [3:0] Pad_Row, Pad_Col,
    output [7:0] row, col
);

    

endmodule